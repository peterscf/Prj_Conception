-----------------------------TOP.vhd----------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;



entity top_num is
   port( 
        i_CLK		   : in  std_logic;                      
	i_RESET_n    	   : in  std_logic;                     
	i_data             : in  std_logic;
	i_in_demod_I	   : in  std_logic_vector(4 downto 0);
	i_in_demod_Q	   : in  std_logic_vector(4 downto 0);
        i_debug_demod      : in  std_logic;
        i_debug_cordic     : in  std_logic;
        o_output           : out std_logic_vector (18 downto 0);
	o_output_comparator: out std_logic_vector (1 downto 0)	
      );
end top_num;

architecture A of top_num is    

------------------------declaration  des composants------------------------------------------
--Modulateur MSK
component msk_modulator is port (	
	i_hclk		: in  std_logic;                      
	i_rstn    : in  std_logic;                     
	i_data    : in  std_logic;   
	o_i       : out std_logic_vector(4 downto 0);  
	o_q       : out std_logic_vector(4 downto 0));  
end component;

--Démodulateur IQ
component Demod_IQ is
  port( 
	I    	    : in  std_logic_vector(4 downto 0);
        Q           : in  std_logic_vector(4 downto 0);
        CLK         : in  std_logic;
        RESET_n     : in  std_logic;
        Filter_outI    : out std_logic_vector(7 downto 0);
        Filter_outQ    : out std_logic_vector(7 downto 0)
      );
end component;

-- CORDIC
component CORDIC_top is
	generic(Nb_b: integer := 8);

	port( 	CLK  : in std_logic;
		RESET_n  : in std_logic;
	  	X  : in  std_logic_vector(Nb_b-1 downto 0);
		Y  : in  std_logic_vector(Nb_b-1 downto 0);
		Z  : out std_logic_vector(8 downto 0));
end component;

component rom_cordic    is 
	port ( 
	CLK      : in std_logic;
	RESET_N  : in std_logic;
	ENABLE   : in std_logic; 
	X        : out std_logic_vector(7 downto 0);
	Y        : out std_logic_vector(7 downto 0)
 	);
end component;


--COMPARATOR
component comparator is 
port(   i_clk       : in std_logic;
	i_restn     : in std_logic;
        i_phase     : in std_logic_vector  (8 downto 0);
        o_comparator: out std_logic_vector (1 downto 0)	
 ); 

end component;
 
------------------------ Fin declaration  des composants------------------------------------------


-- Signaux du Filtre


signal out_modu_I    	: std_logic_vector(4 downto 0);
signal out_modu_Q    	: std_logic_vector(4 downto 0);
signal out_demod_I   	: std_logic_vector(7 downto 0);
signal out_demod_Q   	: std_logic_vector(7 downto 0);   
signal in_cordic_I   	: std_logic_vector(7 downto 0);
signal in_cordic_Q   	: std_logic_vector(7 downto 0);
signal out_phi       	: std_logic_vector(8 downto 0);
signal o_x           	: std_logic_vector(7 downto 0);
signal o_y              : std_logic_vector(7 downto 0);
signal o_out_comparator :  std_logic_vector(1 downto 0);



begin
--Modulateur MSK
modu : msk_modulator  port map (i_CLK, i_RESET_n, i_data, out_modu_I, out_modu_Q);
--Demodulateur IQ
demod : Demod_IQ      port map (i_in_demod_I, i_in_demod_Q, i_CLK, i_RESET_n, out_demod_I, out_demod_Q);
--Cordic
cordic : cordic_top port map (i_CLK, i_RESET_n, in_cordic_I, in_cordic_Q, out_phi);
--Rom_cordic 
rom: rom_cordic   port map (i_CLK,i_RESET_n,i_debug_cordic,o_x,o_y);
--Comparator
comparator_1: comparator port map (i_CLK,i_RESET_n,out_phi,o_out_comparator);


i_cordic_selection:process (i_debug_cordic, out_demod_I, out_demod_Q, o_x, o_y)
begin 
 if (i_debug_cordic = '1' ) then          -- Select Rom
        in_cordic_I <= o_x;
	in_cordic_Q <= o_y; 
 else                                     -- Select Demodulator
	in_cordic_I <= out_demod_I;
	in_cordic_Q <= out_demod_Q;
 end if; 
end process i_cordic_selection;


o_output_selection:process (i_debug_demod, out_demod_I, out_demod_Q, out_modu_I, out_modu_Q, out_phi)
begin
 if (i_debug_demod = '1' ) then          	-- Select Demodulator
 	o_output(18 downto 16) <= "000";
        o_output(15 downto 8) <= out_demod_I;
        o_output(7 downto 0)  <= out_demod_Q; 
 else 						-- Select Cordic and MSK
       o_output(18 downto 14) <= out_modu_I ;
       o_output(13 downto 9) <= out_modu_Q ;
       o_output(8 downto 0) <= out_phi;
 
 end if;

end process o_output_selection;
 

end A;
